// gpu_qsys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module gpu_qsys (
		input  wire        clk_clk,                                 //                               clk.clk
		input  wire [29:0] gpu_main_external_interface_address,     //       gpu_main_external_interface.address
		input  wire [3:0]  gpu_main_external_interface_byte_enable, //                                  .byte_enable
		input  wire        gpu_main_external_interface_read,        //                                  .read
		input  wire        gpu_main_external_interface_write,       //                                  .write
		input  wire [31:0] gpu_main_external_interface_write_data,  //                                  .write_data
		output wire        gpu_main_external_interface_acknowledge, //                                  .acknowledge
		output wire [31:0] gpu_main_external_interface_read_data,   //                                  .read_data
		output wire        instr_fifo_out_valid,                    //                    instr_fifo_out.valid
		output wire [31:0] instr_fifo_out_data,                     //                                  .data
		input  wire        instr_fifo_out_ready,                    //                                  .ready
		output wire [12:0] memory_mem_a,                            //                            memory.mem_a
		output wire [2:0]  memory_mem_ba,                           //                                  .mem_ba
		output wire        memory_mem_ck,                           //                                  .mem_ck
		output wire        memory_mem_ck_n,                         //                                  .mem_ck_n
		output wire        memory_mem_cke,                          //                                  .mem_cke
		output wire        memory_mem_cs_n,                         //                                  .mem_cs_n
		output wire        memory_mem_ras_n,                        //                                  .mem_ras_n
		output wire        memory_mem_cas_n,                        //                                  .mem_cas_n
		output wire        memory_mem_we_n,                         //                                  .mem_we_n
		output wire        memory_mem_reset_n,                      //                                  .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                           //                                  .mem_dq
		inout  wire        memory_mem_dqs,                          //                                  .mem_dqs
		inout  wire        memory_mem_dqs_n,                        //                                  .mem_dqs_n
		output wire        memory_mem_odt,                          //                                  .mem_odt
		output wire        memory_mem_dm,                           //                                  .mem_dm
		input  wire        memory_oct_rzqin,                        //                                  .oct_rzqin
		input  wire        prim_assembly_fifo_in_valid,             //             prim_assembly_fifo_in.valid
		input  wire [31:0] prim_assembly_fifo_in_data,              //                                  .data
		output wire        prim_assembly_fifo_in_ready,             //                                  .ready
		output wire        prim_assembly_fifo_out_valid,            //            prim_assembly_fifo_out.valid
		output wire [31:0] prim_assembly_fifo_out_data,             //                                  .data
		input  wire        prim_assembly_fifo_out_ready,            //                                  .ready
		input  wire        raster_fifo_in_valid,                    //                    raster_fifo_in.valid
		input  wire [31:0] raster_fifo_in_data,                     //                                  .data
		output wire        raster_fifo_in_ready,                    //                                  .ready
		output wire        raster_fifo_out_valid,                   //                   raster_fifo_out.valid
		output wire [31:0] raster_fifo_out_data,                    //                                  .data
		input  wire        raster_fifo_out_ready,                   //                                  .ready
		input  wire        reset_reset,                             //                             reset.reset
		input  wire        vert_processing_fifo_in_valid,           //           vert_processing_fifo_in.valid
		input  wire [31:0] vert_processing_fifo_in_data,            //                                  .data
		output wire        vert_processing_fifo_in_ready,           //                                  .ready
		output wire        vert_processing_fifo_out_valid,          //          vert_processing_fifo_out.valid
		output wire [31:0] vert_processing_fifo_out_data,           //                                  .data
		input  wire        vert_processing_fifo_out_ready,          //                                  .ready
		output wire        vga_controller_external_interface_CLK,   // vga_controller_external_interface.CLK
		output wire        vga_controller_external_interface_HS,    //                                  .HS
		output wire        vga_controller_external_interface_VS,    //                                  .VS
		output wire        vga_controller_external_interface_BLANK, //                                  .BLANK
		output wire        vga_controller_external_interface_SYNC,  //                                  .SYNC
		output wire [7:0]  vga_controller_external_interface_R,     //                                  .R
		output wire [7:0]  vga_controller_external_interface_G,     //                                  .G
		output wire [7:0]  vga_controller_external_interface_B,     //                                  .B
		input  wire        video_pll_ref_clk_clk,                    //                 video_pll_ref_clk.clk
		output wire 			pll_clock,
		output wire				sys_reset
		);

	wire         pixel_fifo_mod_avalon_dc_buffer_source_valid;                         // pixel_fifo_mod:stream_out_valid -> vga_controller:valid
	wire  [29:0] pixel_fifo_mod_avalon_dc_buffer_source_data;                          // pixel_fifo_mod:stream_out_data -> vga_controller:data
	wire         pixel_fifo_mod_avalon_dc_buffer_source_ready;                         // vga_controller:ready -> pixel_fifo_mod:stream_out_ready
	wire         pixel_fifo_mod_avalon_dc_buffer_source_startofpacket;                 // pixel_fifo_mod:stream_out_startofpacket -> vga_controller:startofpacket
	wire         pixel_fifo_mod_avalon_dc_buffer_source_endofpacket;                   // pixel_fifo_mod:stream_out_endofpacket -> vga_controller:endofpacket
	wire         pixel_dma_avalon_pixel_source_valid;                                  // pixel_dma:stream_valid -> pixel_fifo_mod:stream_in_valid
	wire  [29:0] pixel_dma_avalon_pixel_source_data;                                   // pixel_dma:stream_data -> pixel_fifo_mod:stream_in_data
	wire         pixel_dma_avalon_pixel_source_ready;                                  // pixel_fifo_mod:stream_in_ready -> pixel_dma:stream_ready
	wire         pixel_dma_avalon_pixel_source_startofpacket;                          // pixel_dma:stream_startofpacket -> pixel_fifo_mod:stream_in_startofpacket
	wire         pixel_dma_avalon_pixel_source_endofpacket;                            // pixel_dma:stream_endofpacket -> pixel_fifo_mod:stream_in_endofpacket
	wire         pll_outclk0_clk;                                                      // pll:outclk_0 -> [address_span_extender:clk, gpu_main:clk, hps:f2h_axi_clk, hps:f2h_sdram0_clk, hps:h2f_axi_clk, hps:h2f_lw_axi_clk, instr_fifo:rdclock, instr_fifo:wrclock, mm_interconnect_0:pll_outclk0_clk, mm_interconnect_1:pll_outclk0_clk, mm_interconnect_2:pll_outclk0_clk, pixel_dma:clk, pixel_fifo_mod:clk_stream_in, prim_assembly_fifo:rdclock, prim_assembly_fifo:wrclock, raster_fifo:rdclock, raster_fifo:wrclock, rst_controller:clk, vert_processing_fifo:rdclock, vert_processing_fifo:wrclock]
	wire         video_pll_vga_clk_clk;                                                // video_pll:vga_clk_clk -> [pixel_fifo_mod:clk_stream_out, rst_controller_001:clk, vga_controller:clk]
	wire         hps_h2f_reset_reset;                                                  // hps:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0, video_pll:ref_reset_reset]
	wire  [31:0] gpu_main_avalon_master_readdata;                                      // mm_interconnect_0:gpu_main_avalon_master_readdata -> gpu_main:avalon_readdata
	wire         gpu_main_avalon_master_waitrequest;                                   // mm_interconnect_0:gpu_main_avalon_master_waitrequest -> gpu_main:avalon_waitrequest
	wire   [3:0] gpu_main_avalon_master_byteenable;                                    // gpu_main:avalon_byteenable -> mm_interconnect_0:gpu_main_avalon_master_byteenable
	wire         gpu_main_avalon_master_read;                                          // gpu_main:avalon_read -> mm_interconnect_0:gpu_main_avalon_master_read
	wire  [29:0] gpu_main_avalon_master_address;                                       // gpu_main:avalon_address -> mm_interconnect_0:gpu_main_avalon_master_address
	wire         gpu_main_avalon_master_write;                                         // gpu_main:avalon_write -> mm_interconnect_0:gpu_main_avalon_master_write
	wire  [31:0] gpu_main_avalon_master_writedata;                                     // gpu_main:avalon_writedata -> mm_interconnect_0:gpu_main_avalon_master_writedata
	wire  [31:0] mm_interconnect_0_address_span_extender_windowed_slave_readdata;      // address_span_extender:avs_s0_readdata -> mm_interconnect_0:address_span_extender_windowed_slave_readdata
	wire         mm_interconnect_0_address_span_extender_windowed_slave_waitrequest;   // address_span_extender:avs_s0_waitrequest -> mm_interconnect_0:address_span_extender_windowed_slave_waitrequest
	wire  [27:0] mm_interconnect_0_address_span_extender_windowed_slave_address;       // mm_interconnect_0:address_span_extender_windowed_slave_address -> address_span_extender:avs_s0_address
	wire         mm_interconnect_0_address_span_extender_windowed_slave_read;          // mm_interconnect_0:address_span_extender_windowed_slave_read -> address_span_extender:avs_s0_read
	wire   [3:0] mm_interconnect_0_address_span_extender_windowed_slave_byteenable;    // mm_interconnect_0:address_span_extender_windowed_slave_byteenable -> address_span_extender:avs_s0_byteenable
	wire         mm_interconnect_0_address_span_extender_windowed_slave_readdatavalid; // address_span_extender:avs_s0_readdatavalid -> mm_interconnect_0:address_span_extender_windowed_slave_readdatavalid
	wire         mm_interconnect_0_address_span_extender_windowed_slave_write;         // mm_interconnect_0:address_span_extender_windowed_slave_write -> address_span_extender:avs_s0_write
	wire  [31:0] mm_interconnect_0_address_span_extender_windowed_slave_writedata;     // mm_interconnect_0:address_span_extender_windowed_slave_writedata -> address_span_extender:avs_s0_writedata
	wire   [0:0] mm_interconnect_0_address_span_extender_windowed_slave_burstcount;    // mm_interconnect_0:address_span_extender_windowed_slave_burstcount -> address_span_extender:avs_s0_burstcount
	wire         pixel_dma_avalon_pixel_dma_master_waitrequest;                        // mm_interconnect_1:pixel_dma_avalon_pixel_dma_master_waitrequest -> pixel_dma:master_waitrequest
	wire  [31:0] pixel_dma_avalon_pixel_dma_master_readdata;                           // mm_interconnect_1:pixel_dma_avalon_pixel_dma_master_readdata -> pixel_dma:master_readdata
	wire  [31:0] pixel_dma_avalon_pixel_dma_master_address;                            // pixel_dma:master_address -> mm_interconnect_1:pixel_dma_avalon_pixel_dma_master_address
	wire         pixel_dma_avalon_pixel_dma_master_read;                               // pixel_dma:master_read -> mm_interconnect_1:pixel_dma_avalon_pixel_dma_master_read
	wire         pixel_dma_avalon_pixel_dma_master_readdatavalid;                      // mm_interconnect_1:pixel_dma_avalon_pixel_dma_master_readdatavalid -> pixel_dma:master_readdatavalid
	wire         pixel_dma_avalon_pixel_dma_master_lock;                               // pixel_dma:master_arbiterlock -> mm_interconnect_1:pixel_dma_avalon_pixel_dma_master_lock
	wire         address_span_extender_expanded_master_waitrequest;                    // mm_interconnect_1:address_span_extender_expanded_master_waitrequest -> address_span_extender:avm_m0_waitrequest
	wire  [31:0] address_span_extender_expanded_master_readdata;                       // mm_interconnect_1:address_span_extender_expanded_master_readdata -> address_span_extender:avm_m0_readdata
	wire  [31:0] address_span_extender_expanded_master_address;                        // address_span_extender:avm_m0_address -> mm_interconnect_1:address_span_extender_expanded_master_address
	wire         address_span_extender_expanded_master_read;                           // address_span_extender:avm_m0_read -> mm_interconnect_1:address_span_extender_expanded_master_read
	wire   [3:0] address_span_extender_expanded_master_byteenable;                     // address_span_extender:avm_m0_byteenable -> mm_interconnect_1:address_span_extender_expanded_master_byteenable
	wire         address_span_extender_expanded_master_readdatavalid;                  // mm_interconnect_1:address_span_extender_expanded_master_readdatavalid -> address_span_extender:avm_m0_readdatavalid
	wire         address_span_extender_expanded_master_write;                          // address_span_extender:avm_m0_write -> mm_interconnect_1:address_span_extender_expanded_master_write
	wire  [31:0] address_span_extender_expanded_master_writedata;                      // address_span_extender:avm_m0_writedata -> mm_interconnect_1:address_span_extender_expanded_master_writedata
	wire   [0:0] address_span_extender_expanded_master_burstcount;                     // address_span_extender:avm_m0_burstcount -> mm_interconnect_1:address_span_extender_expanded_master_burstcount
	wire   [1:0] mm_interconnect_1_hps_f2h_axi_slave_awburst;                          // mm_interconnect_1:hps_f2h_axi_slave_awburst -> hps:f2h_AWBURST
	wire   [4:0] mm_interconnect_1_hps_f2h_axi_slave_awuser;                           // mm_interconnect_1:hps_f2h_axi_slave_awuser -> hps:f2h_AWUSER
	wire   [3:0] mm_interconnect_1_hps_f2h_axi_slave_arlen;                            // mm_interconnect_1:hps_f2h_axi_slave_arlen -> hps:f2h_ARLEN
	wire   [3:0] mm_interconnect_1_hps_f2h_axi_slave_wstrb;                            // mm_interconnect_1:hps_f2h_axi_slave_wstrb -> hps:f2h_WSTRB
	wire         mm_interconnect_1_hps_f2h_axi_slave_wready;                           // hps:f2h_WREADY -> mm_interconnect_1:hps_f2h_axi_slave_wready
	wire   [7:0] mm_interconnect_1_hps_f2h_axi_slave_rid;                              // hps:f2h_RID -> mm_interconnect_1:hps_f2h_axi_slave_rid
	wire         mm_interconnect_1_hps_f2h_axi_slave_rready;                           // mm_interconnect_1:hps_f2h_axi_slave_rready -> hps:f2h_RREADY
	wire   [3:0] mm_interconnect_1_hps_f2h_axi_slave_awlen;                            // mm_interconnect_1:hps_f2h_axi_slave_awlen -> hps:f2h_AWLEN
	wire   [7:0] mm_interconnect_1_hps_f2h_axi_slave_wid;                              // mm_interconnect_1:hps_f2h_axi_slave_wid -> hps:f2h_WID
	wire   [3:0] mm_interconnect_1_hps_f2h_axi_slave_arcache;                          // mm_interconnect_1:hps_f2h_axi_slave_arcache -> hps:f2h_ARCACHE
	wire         mm_interconnect_1_hps_f2h_axi_slave_wvalid;                           // mm_interconnect_1:hps_f2h_axi_slave_wvalid -> hps:f2h_WVALID
	wire  [31:0] mm_interconnect_1_hps_f2h_axi_slave_araddr;                           // mm_interconnect_1:hps_f2h_axi_slave_araddr -> hps:f2h_ARADDR
	wire   [2:0] mm_interconnect_1_hps_f2h_axi_slave_arprot;                           // mm_interconnect_1:hps_f2h_axi_slave_arprot -> hps:f2h_ARPROT
	wire   [2:0] mm_interconnect_1_hps_f2h_axi_slave_awprot;                           // mm_interconnect_1:hps_f2h_axi_slave_awprot -> hps:f2h_AWPROT
	wire  [31:0] mm_interconnect_1_hps_f2h_axi_slave_wdata;                            // mm_interconnect_1:hps_f2h_axi_slave_wdata -> hps:f2h_WDATA
	wire         mm_interconnect_1_hps_f2h_axi_slave_arvalid;                          // mm_interconnect_1:hps_f2h_axi_slave_arvalid -> hps:f2h_ARVALID
	wire   [3:0] mm_interconnect_1_hps_f2h_axi_slave_awcache;                          // mm_interconnect_1:hps_f2h_axi_slave_awcache -> hps:f2h_AWCACHE
	wire   [7:0] mm_interconnect_1_hps_f2h_axi_slave_arid;                             // mm_interconnect_1:hps_f2h_axi_slave_arid -> hps:f2h_ARID
	wire   [1:0] mm_interconnect_1_hps_f2h_axi_slave_arlock;                           // mm_interconnect_1:hps_f2h_axi_slave_arlock -> hps:f2h_ARLOCK
	wire   [1:0] mm_interconnect_1_hps_f2h_axi_slave_awlock;                           // mm_interconnect_1:hps_f2h_axi_slave_awlock -> hps:f2h_AWLOCK
	wire  [31:0] mm_interconnect_1_hps_f2h_axi_slave_awaddr;                           // mm_interconnect_1:hps_f2h_axi_slave_awaddr -> hps:f2h_AWADDR
	wire   [1:0] mm_interconnect_1_hps_f2h_axi_slave_bresp;                            // hps:f2h_BRESP -> mm_interconnect_1:hps_f2h_axi_slave_bresp
	wire         mm_interconnect_1_hps_f2h_axi_slave_arready;                          // hps:f2h_ARREADY -> mm_interconnect_1:hps_f2h_axi_slave_arready
	wire  [31:0] mm_interconnect_1_hps_f2h_axi_slave_rdata;                            // hps:f2h_RDATA -> mm_interconnect_1:hps_f2h_axi_slave_rdata
	wire         mm_interconnect_1_hps_f2h_axi_slave_awready;                          // hps:f2h_AWREADY -> mm_interconnect_1:hps_f2h_axi_slave_awready
	wire   [1:0] mm_interconnect_1_hps_f2h_axi_slave_arburst;                          // mm_interconnect_1:hps_f2h_axi_slave_arburst -> hps:f2h_ARBURST
	wire   [2:0] mm_interconnect_1_hps_f2h_axi_slave_arsize;                           // mm_interconnect_1:hps_f2h_axi_slave_arsize -> hps:f2h_ARSIZE
	wire         mm_interconnect_1_hps_f2h_axi_slave_bready;                           // mm_interconnect_1:hps_f2h_axi_slave_bready -> hps:f2h_BREADY
	wire         mm_interconnect_1_hps_f2h_axi_slave_rlast;                            // hps:f2h_RLAST -> mm_interconnect_1:hps_f2h_axi_slave_rlast
	wire         mm_interconnect_1_hps_f2h_axi_slave_wlast;                            // mm_interconnect_1:hps_f2h_axi_slave_wlast -> hps:f2h_WLAST
	wire   [1:0] mm_interconnect_1_hps_f2h_axi_slave_rresp;                            // hps:f2h_RRESP -> mm_interconnect_1:hps_f2h_axi_slave_rresp
	wire   [7:0] mm_interconnect_1_hps_f2h_axi_slave_awid;                             // mm_interconnect_1:hps_f2h_axi_slave_awid -> hps:f2h_AWID
	wire   [7:0] mm_interconnect_1_hps_f2h_axi_slave_bid;                              // hps:f2h_BID -> mm_interconnect_1:hps_f2h_axi_slave_bid
	wire         mm_interconnect_1_hps_f2h_axi_slave_bvalid;                           // hps:f2h_BVALID -> mm_interconnect_1:hps_f2h_axi_slave_bvalid
	wire   [2:0] mm_interconnect_1_hps_f2h_axi_slave_awsize;                           // mm_interconnect_1:hps_f2h_axi_slave_awsize -> hps:f2h_AWSIZE
	wire         mm_interconnect_1_hps_f2h_axi_slave_awvalid;                          // mm_interconnect_1:hps_f2h_axi_slave_awvalid -> hps:f2h_AWVALID
	wire   [4:0] mm_interconnect_1_hps_f2h_axi_slave_aruser;                           // mm_interconnect_1:hps_f2h_axi_slave_aruser -> hps:f2h_ARUSER
	wire         mm_interconnect_1_hps_f2h_axi_slave_rvalid;                           // hps:f2h_RVALID -> mm_interconnect_1:hps_f2h_axi_slave_rvalid
	wire   [1:0] hps_h2f_axi_master_awburst;                                           // hps:h2f_AWBURST -> mm_interconnect_2:hps_h2f_axi_master_awburst
	wire   [3:0] hps_h2f_axi_master_arlen;                                             // hps:h2f_ARLEN -> mm_interconnect_2:hps_h2f_axi_master_arlen
	wire   [3:0] hps_h2f_axi_master_wstrb;                                             // hps:h2f_WSTRB -> mm_interconnect_2:hps_h2f_axi_master_wstrb
	wire         hps_h2f_axi_master_wready;                                            // mm_interconnect_2:hps_h2f_axi_master_wready -> hps:h2f_WREADY
	wire  [11:0] hps_h2f_axi_master_rid;                                               // mm_interconnect_2:hps_h2f_axi_master_rid -> hps:h2f_RID
	wire         hps_h2f_axi_master_rready;                                            // hps:h2f_RREADY -> mm_interconnect_2:hps_h2f_axi_master_rready
	wire   [3:0] hps_h2f_axi_master_awlen;                                             // hps:h2f_AWLEN -> mm_interconnect_2:hps_h2f_axi_master_awlen
	wire  [11:0] hps_h2f_axi_master_wid;                                               // hps:h2f_WID -> mm_interconnect_2:hps_h2f_axi_master_wid
	wire   [3:0] hps_h2f_axi_master_arcache;                                           // hps:h2f_ARCACHE -> mm_interconnect_2:hps_h2f_axi_master_arcache
	wire         hps_h2f_axi_master_wvalid;                                            // hps:h2f_WVALID -> mm_interconnect_2:hps_h2f_axi_master_wvalid
	wire  [29:0] hps_h2f_axi_master_araddr;                                            // hps:h2f_ARADDR -> mm_interconnect_2:hps_h2f_axi_master_araddr
	wire   [2:0] hps_h2f_axi_master_arprot;                                            // hps:h2f_ARPROT -> mm_interconnect_2:hps_h2f_axi_master_arprot
	wire   [2:0] hps_h2f_axi_master_awprot;                                            // hps:h2f_AWPROT -> mm_interconnect_2:hps_h2f_axi_master_awprot
	wire  [31:0] hps_h2f_axi_master_wdata;                                             // hps:h2f_WDATA -> mm_interconnect_2:hps_h2f_axi_master_wdata
	wire         hps_h2f_axi_master_arvalid;                                           // hps:h2f_ARVALID -> mm_interconnect_2:hps_h2f_axi_master_arvalid
	wire   [3:0] hps_h2f_axi_master_awcache;                                           // hps:h2f_AWCACHE -> mm_interconnect_2:hps_h2f_axi_master_awcache
	wire  [11:0] hps_h2f_axi_master_arid;                                              // hps:h2f_ARID -> mm_interconnect_2:hps_h2f_axi_master_arid
	wire   [1:0] hps_h2f_axi_master_arlock;                                            // hps:h2f_ARLOCK -> mm_interconnect_2:hps_h2f_axi_master_arlock
	wire   [1:0] hps_h2f_axi_master_awlock;                                            // hps:h2f_AWLOCK -> mm_interconnect_2:hps_h2f_axi_master_awlock
	wire  [29:0] hps_h2f_axi_master_awaddr;                                            // hps:h2f_AWADDR -> mm_interconnect_2:hps_h2f_axi_master_awaddr
	wire   [1:0] hps_h2f_axi_master_bresp;                                             // mm_interconnect_2:hps_h2f_axi_master_bresp -> hps:h2f_BRESP
	wire         hps_h2f_axi_master_arready;                                           // mm_interconnect_2:hps_h2f_axi_master_arready -> hps:h2f_ARREADY
	wire  [31:0] hps_h2f_axi_master_rdata;                                             // mm_interconnect_2:hps_h2f_axi_master_rdata -> hps:h2f_RDATA
	wire         hps_h2f_axi_master_awready;                                           // mm_interconnect_2:hps_h2f_axi_master_awready -> hps:h2f_AWREADY
	wire   [1:0] hps_h2f_axi_master_arburst;                                           // hps:h2f_ARBURST -> mm_interconnect_2:hps_h2f_axi_master_arburst
	wire   [2:0] hps_h2f_axi_master_arsize;                                            // hps:h2f_ARSIZE -> mm_interconnect_2:hps_h2f_axi_master_arsize
	wire         hps_h2f_axi_master_bready;                                            // hps:h2f_BREADY -> mm_interconnect_2:hps_h2f_axi_master_bready
	wire         hps_h2f_axi_master_rlast;                                             // mm_interconnect_2:hps_h2f_axi_master_rlast -> hps:h2f_RLAST
	wire         hps_h2f_axi_master_wlast;                                             // hps:h2f_WLAST -> mm_interconnect_2:hps_h2f_axi_master_wlast
	wire   [1:0] hps_h2f_axi_master_rresp;                                             // mm_interconnect_2:hps_h2f_axi_master_rresp -> hps:h2f_RRESP
	wire  [11:0] hps_h2f_axi_master_awid;                                              // hps:h2f_AWID -> mm_interconnect_2:hps_h2f_axi_master_awid
	wire  [11:0] hps_h2f_axi_master_bid;                                               // mm_interconnect_2:hps_h2f_axi_master_bid -> hps:h2f_BID
	wire         hps_h2f_axi_master_bvalid;                                            // mm_interconnect_2:hps_h2f_axi_master_bvalid -> hps:h2f_BVALID
	wire   [2:0] hps_h2f_axi_master_awsize;                                            // hps:h2f_AWSIZE -> mm_interconnect_2:hps_h2f_axi_master_awsize
	wire         hps_h2f_axi_master_awvalid;                                           // hps:h2f_AWVALID -> mm_interconnect_2:hps_h2f_axi_master_awvalid
	wire         hps_h2f_axi_master_rvalid;                                            // mm_interconnect_2:hps_h2f_axi_master_rvalid -> hps:h2f_RVALID
	wire  [31:0] mm_interconnect_2_pixel_dma_avalon_control_slave_readdata;            // pixel_dma:slave_readdata -> mm_interconnect_2:pixel_dma_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_2_pixel_dma_avalon_control_slave_address;             // mm_interconnect_2:pixel_dma_avalon_control_slave_address -> pixel_dma:slave_address
	wire         mm_interconnect_2_pixel_dma_avalon_control_slave_read;                // mm_interconnect_2:pixel_dma_avalon_control_slave_read -> pixel_dma:slave_read
	wire   [3:0] mm_interconnect_2_pixel_dma_avalon_control_slave_byteenable;          // mm_interconnect_2:pixel_dma_avalon_control_slave_byteenable -> pixel_dma:slave_byteenable
	wire         mm_interconnect_2_pixel_dma_avalon_control_slave_write;               // mm_interconnect_2:pixel_dma_avalon_control_slave_write -> pixel_dma:slave_write
	wire  [31:0] mm_interconnect_2_pixel_dma_avalon_control_slave_writedata;           // mm_interconnect_2:pixel_dma_avalon_control_slave_writedata -> pixel_dma:slave_writedata
	wire         mm_interconnect_2_instr_fifo_in_waitrequest;                          // instr_fifo:avalonmm_write_slave_waitrequest -> mm_interconnect_2:instr_fifo_in_waitrequest
	wire   [0:0] mm_interconnect_2_instr_fifo_in_address;                              // mm_interconnect_2:instr_fifo_in_address -> instr_fifo:avalonmm_write_slave_address
	wire         mm_interconnect_2_instr_fifo_in_write;                                // mm_interconnect_2:instr_fifo_in_write -> instr_fifo:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_2_instr_fifo_in_writedata;                            // mm_interconnect_2:instr_fifo_in_writedata -> instr_fifo:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_2_instr_fifo_in_csr_readdata;                         // instr_fifo:wrclk_control_slave_readdata -> mm_interconnect_2:instr_fifo_in_csr_readdata
	wire   [2:0] mm_interconnect_2_instr_fifo_in_csr_address;                          // mm_interconnect_2:instr_fifo_in_csr_address -> instr_fifo:wrclk_control_slave_address
	wire         mm_interconnect_2_instr_fifo_in_csr_read;                             // mm_interconnect_2:instr_fifo_in_csr_read -> instr_fifo:wrclk_control_slave_read
	wire         mm_interconnect_2_instr_fifo_in_csr_write;                            // mm_interconnect_2:instr_fifo_in_csr_write -> instr_fifo:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_2_instr_fifo_in_csr_writedata;                        // mm_interconnect_2:instr_fifo_in_csr_writedata -> instr_fifo:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_2_vert_processing_fifo_out_csr_readdata;              // vert_processing_fifo:rdclk_control_slave_readdata -> mm_interconnect_2:vert_processing_fifo_out_csr_readdata
	wire   [2:0] mm_interconnect_2_vert_processing_fifo_out_csr_address;               // mm_interconnect_2:vert_processing_fifo_out_csr_address -> vert_processing_fifo:rdclk_control_slave_address
	wire         mm_interconnect_2_vert_processing_fifo_out_csr_read;                  // mm_interconnect_2:vert_processing_fifo_out_csr_read -> vert_processing_fifo:rdclk_control_slave_read
	wire         mm_interconnect_2_vert_processing_fifo_out_csr_write;                 // mm_interconnect_2:vert_processing_fifo_out_csr_write -> vert_processing_fifo:rdclk_control_slave_write
	wire  [31:0] mm_interconnect_2_vert_processing_fifo_out_csr_writedata;             // mm_interconnect_2:vert_processing_fifo_out_csr_writedata -> vert_processing_fifo:rdclk_control_slave_writedata
	wire  [31:0] mm_interconnect_2_prim_assembly_fifo_out_csr_readdata;                // prim_assembly_fifo:rdclk_control_slave_readdata -> mm_interconnect_2:prim_assembly_fifo_out_csr_readdata
	wire   [2:0] mm_interconnect_2_prim_assembly_fifo_out_csr_address;                 // mm_interconnect_2:prim_assembly_fifo_out_csr_address -> prim_assembly_fifo:rdclk_control_slave_address
	wire         mm_interconnect_2_prim_assembly_fifo_out_csr_read;                    // mm_interconnect_2:prim_assembly_fifo_out_csr_read -> prim_assembly_fifo:rdclk_control_slave_read
	wire         mm_interconnect_2_prim_assembly_fifo_out_csr_write;                   // mm_interconnect_2:prim_assembly_fifo_out_csr_write -> prim_assembly_fifo:rdclk_control_slave_write
	wire  [31:0] mm_interconnect_2_prim_assembly_fifo_out_csr_writedata;               // mm_interconnect_2:prim_assembly_fifo_out_csr_writedata -> prim_assembly_fifo:rdclk_control_slave_writedata
	wire  [31:0] mm_interconnect_2_raster_fifo_out_csr_readdata;                       // raster_fifo:rdclk_control_slave_readdata -> mm_interconnect_2:raster_fifo_out_csr_readdata
	wire   [2:0] mm_interconnect_2_raster_fifo_out_csr_address;                        // mm_interconnect_2:raster_fifo_out_csr_address -> raster_fifo:rdclk_control_slave_address
	wire         mm_interconnect_2_raster_fifo_out_csr_read;                           // mm_interconnect_2:raster_fifo_out_csr_read -> raster_fifo:rdclk_control_slave_read
	wire         mm_interconnect_2_raster_fifo_out_csr_write;                          // mm_interconnect_2:raster_fifo_out_csr_write -> raster_fifo:rdclk_control_slave_write
	wire  [31:0] mm_interconnect_2_raster_fifo_out_csr_writedata;                      // mm_interconnect_2:raster_fifo_out_csr_writedata -> raster_fifo:rdclk_control_slave_writedata
	wire         rst_controller_reset_out_reset;                                       // rst_controller:reset_out -> [address_span_extender:reset, gpu_main:reset, instr_fifo:rdreset_n, instr_fifo:wrreset_n, mm_interconnect_0:gpu_main_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pixel_dma_reset_reset_bridge_in_reset_reset, mm_interconnect_2:pixel_dma_reset_reset_bridge_in_reset_reset, pixel_dma:reset, pixel_fifo_mod:reset_stream_in, prim_assembly_fifo:rdreset_n, prim_assembly_fifo:wrreset_n, raster_fifo:rdreset_n, raster_fifo:wrreset_n, vert_processing_fifo:rdreset_n, vert_processing_fifo:wrreset_n]
	wire         rst_controller_001_reset_out_reset;                                   // rst_controller_001:reset_out -> [pixel_fifo_mod:reset_stream_out, vga_controller:reset]
	wire         video_pll_reset_source_reset;                                         // video_pll:reset_source_reset -> rst_controller_001:reset_in1

	assign sys_reset = rst_controller_reset_out_reset;
	assign pll_clock = pll_outclk0_clk;
	
	altera_address_span_extender #(
		.DATA_WIDTH           (32),
		.BYTEENABLE_WIDTH     (4),
		.MASTER_ADDRESS_WIDTH (32),
		.SLAVE_ADDRESS_WIDTH  (28),
		.SLAVE_ADDRESS_SHIFT  (2),
		.BURSTCOUNT_WIDTH     (1),
		.CNTL_ADDRESS_WIDTH   (1),
		.SUB_WINDOW_COUNT     (1),
		.MASTER_ADDRESS_DEF   (64'b0000000000000000000000000000000000000000000000000000000000000000)
	) address_span_extender (
		.clk                  (pll_outclk0_clk),                                                      //           clock.clk
		.reset                (rst_controller_reset_out_reset),                                       //           reset.reset
		.avs_s0_address       (mm_interconnect_0_address_span_extender_windowed_slave_address),       //  windowed_slave.address
		.avs_s0_read          (mm_interconnect_0_address_span_extender_windowed_slave_read),          //                .read
		.avs_s0_readdata      (mm_interconnect_0_address_span_extender_windowed_slave_readdata),      //                .readdata
		.avs_s0_write         (mm_interconnect_0_address_span_extender_windowed_slave_write),         //                .write
		.avs_s0_writedata     (mm_interconnect_0_address_span_extender_windowed_slave_writedata),     //                .writedata
		.avs_s0_readdatavalid (mm_interconnect_0_address_span_extender_windowed_slave_readdatavalid), //                .readdatavalid
		.avs_s0_waitrequest   (mm_interconnect_0_address_span_extender_windowed_slave_waitrequest),   //                .waitrequest
		.avs_s0_byteenable    (mm_interconnect_0_address_span_extender_windowed_slave_byteenable),    //                .byteenable
		.avs_s0_burstcount    (mm_interconnect_0_address_span_extender_windowed_slave_burstcount),    //                .burstcount
		.avm_m0_address       (address_span_extender_expanded_master_address),                        // expanded_master.address
		.avm_m0_read          (address_span_extender_expanded_master_read),                           //                .read
		.avm_m0_waitrequest   (address_span_extender_expanded_master_waitrequest),                    //                .waitrequest
		.avm_m0_readdata      (address_span_extender_expanded_master_readdata),                       //                .readdata
		.avm_m0_write         (address_span_extender_expanded_master_write),                          //                .write
		.avm_m0_writedata     (address_span_extender_expanded_master_writedata),                      //                .writedata
		.avm_m0_readdatavalid (address_span_extender_expanded_master_readdatavalid),                  //                .readdatavalid
		.avm_m0_byteenable    (address_span_extender_expanded_master_byteenable),                     //                .byteenable
		.avm_m0_burstcount    (address_span_extender_expanded_master_burstcount),                     //                .burstcount
		.avs_cntl_address     (1'b0),                                                                 //     (terminated)
		.avs_cntl_read        (1'b0),                                                                 //     (terminated)
		.avs_cntl_readdata    (),                                                                     //     (terminated)
		.avs_cntl_write       (1'b0),                                                                 //     (terminated)
		.avs_cntl_writedata   (64'b0000000000000000000000000000000000000000000000000000000000000000), //     (terminated)
		.avs_cntl_byteenable  (8'b00000000)                                                           //     (terminated)
	);

	gpu_qsys_gpu_main gpu_main (
		.clk                (pll_outclk0_clk),                         //                clk.clk
		.reset              (rst_controller_reset_out_reset),          //              reset.reset
		.avalon_readdata    (gpu_main_avalon_master_readdata),         //      avalon_master.readdata
		.avalon_waitrequest (gpu_main_avalon_master_waitrequest),      //                   .waitrequest
		.avalon_byteenable  (gpu_main_avalon_master_byteenable),       //                   .byteenable
		.avalon_read        (gpu_main_avalon_master_read),             //                   .read
		.avalon_write       (gpu_main_avalon_master_write),            //                   .write
		.avalon_writedata   (gpu_main_avalon_master_writedata),        //                   .writedata
		.avalon_address     (gpu_main_avalon_master_address),          //                   .address
		.address            (gpu_main_external_interface_address),     // external_interface.export
		.byte_enable        (gpu_main_external_interface_byte_enable), //                   .export
		.read               (gpu_main_external_interface_read),        //                   .export
		.write              (gpu_main_external_interface_write),       //                   .export
		.write_data         (gpu_main_external_interface_write_data),  //                   .export
		.acknowledge        (gpu_main_external_interface_acknowledge), //                   .export
		.read_data          (gpu_main_external_interface_read_data)    //                   .export
	);

	gpu_qsys_hps #(
		.F2S_Width (1),
		.S2F_Width (1)
	) hps (
		.mem_a                  (memory_mem_a),                                //            memory.mem_a
		.mem_ba                 (memory_mem_ba),                               //                  .mem_ba
		.mem_ck                 (memory_mem_ck),                               //                  .mem_ck
		.mem_ck_n               (memory_mem_ck_n),                             //                  .mem_ck_n
		.mem_cke                (memory_mem_cke),                              //                  .mem_cke
		.mem_cs_n               (memory_mem_cs_n),                             //                  .mem_cs_n
		.mem_ras_n              (memory_mem_ras_n),                            //                  .mem_ras_n
		.mem_cas_n              (memory_mem_cas_n),                            //                  .mem_cas_n
		.mem_we_n               (memory_mem_we_n),                             //                  .mem_we_n
		.mem_reset_n            (memory_mem_reset_n),                          //                  .mem_reset_n
		.mem_dq                 (memory_mem_dq),                               //                  .mem_dq
		.mem_dqs                (memory_mem_dqs),                              //                  .mem_dqs
		.mem_dqs_n              (memory_mem_dqs_n),                            //                  .mem_dqs_n
		.mem_odt                (memory_mem_odt),                              //                  .mem_odt
		.mem_dm                 (memory_mem_dm),                               //                  .mem_dm
		.oct_rzqin              (memory_oct_rzqin),                            //                  .oct_rzqin
		.h2f_rst_n              (hps_h2f_reset_reset),                         //         h2f_reset.reset_n
		.f2h_sdram0_clk         (pll_outclk0_clk),                             //  f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS     (),                                            //   f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT  (),                                            //                  .burstcount
		.f2h_sdram0_WAITREQUEST (),                                            //                  .waitrequest
		.f2h_sdram0_WRITEDATA   (),                                            //                  .writedata
		.f2h_sdram0_BYTEENABLE  (),                                            //                  .byteenable
		.f2h_sdram0_WRITE       (),                                            //                  .write
		.h2f_axi_clk            (pll_outclk0_clk),                             //     h2f_axi_clock.clk
		.h2f_AWID               (hps_h2f_axi_master_awid),                     //    h2f_axi_master.awid
		.h2f_AWADDR             (hps_h2f_axi_master_awaddr),                   //                  .awaddr
		.h2f_AWLEN              (hps_h2f_axi_master_awlen),                    //                  .awlen
		.h2f_AWSIZE             (hps_h2f_axi_master_awsize),                   //                  .awsize
		.h2f_AWBURST            (hps_h2f_axi_master_awburst),                  //                  .awburst
		.h2f_AWLOCK             (hps_h2f_axi_master_awlock),                   //                  .awlock
		.h2f_AWCACHE            (hps_h2f_axi_master_awcache),                  //                  .awcache
		.h2f_AWPROT             (hps_h2f_axi_master_awprot),                   //                  .awprot
		.h2f_AWVALID            (hps_h2f_axi_master_awvalid),                  //                  .awvalid
		.h2f_AWREADY            (hps_h2f_axi_master_awready),                  //                  .awready
		.h2f_WID                (hps_h2f_axi_master_wid),                      //                  .wid
		.h2f_WDATA              (hps_h2f_axi_master_wdata),                    //                  .wdata
		.h2f_WSTRB              (hps_h2f_axi_master_wstrb),                    //                  .wstrb
		.h2f_WLAST              (hps_h2f_axi_master_wlast),                    //                  .wlast
		.h2f_WVALID             (hps_h2f_axi_master_wvalid),                   //                  .wvalid
		.h2f_WREADY             (hps_h2f_axi_master_wready),                   //                  .wready
		.h2f_BID                (hps_h2f_axi_master_bid),                      //                  .bid
		.h2f_BRESP              (hps_h2f_axi_master_bresp),                    //                  .bresp
		.h2f_BVALID             (hps_h2f_axi_master_bvalid),                   //                  .bvalid
		.h2f_BREADY             (hps_h2f_axi_master_bready),                   //                  .bready
		.h2f_ARID               (hps_h2f_axi_master_arid),                     //                  .arid
		.h2f_ARADDR             (hps_h2f_axi_master_araddr),                   //                  .araddr
		.h2f_ARLEN              (hps_h2f_axi_master_arlen),                    //                  .arlen
		.h2f_ARSIZE             (hps_h2f_axi_master_arsize),                   //                  .arsize
		.h2f_ARBURST            (hps_h2f_axi_master_arburst),                  //                  .arburst
		.h2f_ARLOCK             (hps_h2f_axi_master_arlock),                   //                  .arlock
		.h2f_ARCACHE            (hps_h2f_axi_master_arcache),                  //                  .arcache
		.h2f_ARPROT             (hps_h2f_axi_master_arprot),                   //                  .arprot
		.h2f_ARVALID            (hps_h2f_axi_master_arvalid),                  //                  .arvalid
		.h2f_ARREADY            (hps_h2f_axi_master_arready),                  //                  .arready
		.h2f_RID                (hps_h2f_axi_master_rid),                      //                  .rid
		.h2f_RDATA              (hps_h2f_axi_master_rdata),                    //                  .rdata
		.h2f_RRESP              (hps_h2f_axi_master_rresp),                    //                  .rresp
		.h2f_RLAST              (hps_h2f_axi_master_rlast),                    //                  .rlast
		.h2f_RVALID             (hps_h2f_axi_master_rvalid),                   //                  .rvalid
		.h2f_RREADY             (hps_h2f_axi_master_rready),                   //                  .rready
		.f2h_axi_clk            (pll_outclk0_clk),                             //     f2h_axi_clock.clk
		.f2h_AWID               (mm_interconnect_1_hps_f2h_axi_slave_awid),    //     f2h_axi_slave.awid
		.f2h_AWADDR             (mm_interconnect_1_hps_f2h_axi_slave_awaddr),  //                  .awaddr
		.f2h_AWLEN              (mm_interconnect_1_hps_f2h_axi_slave_awlen),   //                  .awlen
		.f2h_AWSIZE             (mm_interconnect_1_hps_f2h_axi_slave_awsize),  //                  .awsize
		.f2h_AWBURST            (mm_interconnect_1_hps_f2h_axi_slave_awburst), //                  .awburst
		.f2h_AWLOCK             (mm_interconnect_1_hps_f2h_axi_slave_awlock),  //                  .awlock
		.f2h_AWCACHE            (mm_interconnect_1_hps_f2h_axi_slave_awcache), //                  .awcache
		.f2h_AWPROT             (mm_interconnect_1_hps_f2h_axi_slave_awprot),  //                  .awprot
		.f2h_AWVALID            (mm_interconnect_1_hps_f2h_axi_slave_awvalid), //                  .awvalid
		.f2h_AWREADY            (mm_interconnect_1_hps_f2h_axi_slave_awready), //                  .awready
		.f2h_AWUSER             (mm_interconnect_1_hps_f2h_axi_slave_awuser),  //                  .awuser
		.f2h_WID                (mm_interconnect_1_hps_f2h_axi_slave_wid),     //                  .wid
		.f2h_WDATA              (mm_interconnect_1_hps_f2h_axi_slave_wdata),   //                  .wdata
		.f2h_WSTRB              (mm_interconnect_1_hps_f2h_axi_slave_wstrb),   //                  .wstrb
		.f2h_WLAST              (mm_interconnect_1_hps_f2h_axi_slave_wlast),   //                  .wlast
		.f2h_WVALID             (mm_interconnect_1_hps_f2h_axi_slave_wvalid),  //                  .wvalid
		.f2h_WREADY             (mm_interconnect_1_hps_f2h_axi_slave_wready),  //                  .wready
		.f2h_BID                (mm_interconnect_1_hps_f2h_axi_slave_bid),     //                  .bid
		.f2h_BRESP              (mm_interconnect_1_hps_f2h_axi_slave_bresp),   //                  .bresp
		.f2h_BVALID             (mm_interconnect_1_hps_f2h_axi_slave_bvalid),  //                  .bvalid
		.f2h_BREADY             (mm_interconnect_1_hps_f2h_axi_slave_bready),  //                  .bready
		.f2h_ARID               (mm_interconnect_1_hps_f2h_axi_slave_arid),    //                  .arid
		.f2h_ARADDR             (mm_interconnect_1_hps_f2h_axi_slave_araddr),  //                  .araddr
		.f2h_ARLEN              (mm_interconnect_1_hps_f2h_axi_slave_arlen),   //                  .arlen
		.f2h_ARSIZE             (mm_interconnect_1_hps_f2h_axi_slave_arsize),  //                  .arsize
		.f2h_ARBURST            (mm_interconnect_1_hps_f2h_axi_slave_arburst), //                  .arburst
		.f2h_ARLOCK             (mm_interconnect_1_hps_f2h_axi_slave_arlock),  //                  .arlock
		.f2h_ARCACHE            (mm_interconnect_1_hps_f2h_axi_slave_arcache), //                  .arcache
		.f2h_ARPROT             (mm_interconnect_1_hps_f2h_axi_slave_arprot),  //                  .arprot
		.f2h_ARVALID            (mm_interconnect_1_hps_f2h_axi_slave_arvalid), //                  .arvalid
		.f2h_ARREADY            (mm_interconnect_1_hps_f2h_axi_slave_arready), //                  .arready
		.f2h_ARUSER             (mm_interconnect_1_hps_f2h_axi_slave_aruser),  //                  .aruser
		.f2h_RID                (mm_interconnect_1_hps_f2h_axi_slave_rid),     //                  .rid
		.f2h_RDATA              (mm_interconnect_1_hps_f2h_axi_slave_rdata),   //                  .rdata
		.f2h_RRESP              (mm_interconnect_1_hps_f2h_axi_slave_rresp),   //                  .rresp
		.f2h_RLAST              (mm_interconnect_1_hps_f2h_axi_slave_rlast),   //                  .rlast
		.f2h_RVALID             (mm_interconnect_1_hps_f2h_axi_slave_rvalid),  //                  .rvalid
		.f2h_RREADY             (mm_interconnect_1_hps_f2h_axi_slave_rready),  //                  .rready
		.h2f_lw_axi_clk         (pll_outclk0_clk),                             //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID            (),                                            // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR          (),                                            //                  .awaddr
		.h2f_lw_AWLEN           (),                                            //                  .awlen
		.h2f_lw_AWSIZE          (),                                            //                  .awsize
		.h2f_lw_AWBURST         (),                                            //                  .awburst
		.h2f_lw_AWLOCK          (),                                            //                  .awlock
		.h2f_lw_AWCACHE         (),                                            //                  .awcache
		.h2f_lw_AWPROT          (),                                            //                  .awprot
		.h2f_lw_AWVALID         (),                                            //                  .awvalid
		.h2f_lw_AWREADY         (),                                            //                  .awready
		.h2f_lw_WID             (),                                            //                  .wid
		.h2f_lw_WDATA           (),                                            //                  .wdata
		.h2f_lw_WSTRB           (),                                            //                  .wstrb
		.h2f_lw_WLAST           (),                                            //                  .wlast
		.h2f_lw_WVALID          (),                                            //                  .wvalid
		.h2f_lw_WREADY          (),                                            //                  .wready
		.h2f_lw_BID             (),                                            //                  .bid
		.h2f_lw_BRESP           (),                                            //                  .bresp
		.h2f_lw_BVALID          (),                                            //                  .bvalid
		.h2f_lw_BREADY          (),                                            //                  .bready
		.h2f_lw_ARID            (),                                            //                  .arid
		.h2f_lw_ARADDR          (),                                            //                  .araddr
		.h2f_lw_ARLEN           (),                                            //                  .arlen
		.h2f_lw_ARSIZE          (),                                            //                  .arsize
		.h2f_lw_ARBURST         (),                                            //                  .arburst
		.h2f_lw_ARLOCK          (),                                            //                  .arlock
		.h2f_lw_ARCACHE         (),                                            //                  .arcache
		.h2f_lw_ARPROT          (),                                            //                  .arprot
		.h2f_lw_ARVALID         (),                                            //                  .arvalid
		.h2f_lw_ARREADY         (),                                            //                  .arready
		.h2f_lw_RID             (),                                            //                  .rid
		.h2f_lw_RDATA           (),                                            //                  .rdata
		.h2f_lw_RRESP           (),                                            //                  .rresp
		.h2f_lw_RLAST           (),                                            //                  .rlast
		.h2f_lw_RVALID          (),                                            //                  .rvalid
		.h2f_lw_RREADY          ()                                             //                  .rready
	);

	gpu_qsys_instr_fifo instr_fifo (
		.wrclock                          (pll_outclk0_clk),                               //    clk_in.clk
		.wrreset_n                        (~rst_controller_reset_out_reset),               //  reset_in.reset_n
		.rdclock                          (pll_outclk0_clk),                               //   clk_out.clk
		.rdreset_n                        (~rst_controller_reset_out_reset),               // reset_out.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_2_instr_fifo_in_writedata),     //        in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_2_instr_fifo_in_write),         //          .write
		.avalonmm_write_slave_address     (mm_interconnect_2_instr_fifo_in_address),       //          .address
		.avalonmm_write_slave_waitrequest (mm_interconnect_2_instr_fifo_in_waitrequest),   //          .waitrequest
		.avalonst_source_valid            (instr_fifo_out_valid),                          //       out.valid
		.avalonst_source_data             (instr_fifo_out_data),                           //          .data
		.avalonst_source_ready            (instr_fifo_out_ready),                          //          .ready
		.rdclk_control_slave_address      (),                                              //   out_csr.address
		.rdclk_control_slave_read         (),                                              //          .read
		.rdclk_control_slave_writedata    (),                                              //          .writedata
		.rdclk_control_slave_write        (),                                              //          .write
		.rdclk_control_slave_readdata     (),                                              //          .readdata
		.wrclk_control_slave_address      (mm_interconnect_2_instr_fifo_in_csr_address),   //    in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_2_instr_fifo_in_csr_read),      //          .read
		.wrclk_control_slave_writedata    (mm_interconnect_2_instr_fifo_in_csr_writedata), //          .writedata
		.wrclk_control_slave_write        (mm_interconnect_2_instr_fifo_in_csr_write),     //          .write
		.wrclk_control_slave_readdata     (mm_interconnect_2_instr_fifo_in_csr_readdata)   //          .readdata
	);

	gpu_qsys_pixel_dma pixel_dma (
		.clk                  (pll_outclk0_clk),                                             //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                              //                   reset.reset
		.master_readdatavalid (pixel_dma_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_dma_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (pixel_dma_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (pixel_dma_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (pixel_dma_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (pixel_dma_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_2_pixel_dma_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_2_pixel_dma_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_2_pixel_dma_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_2_pixel_dma_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_2_pixel_dma_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_2_pixel_dma_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (pixel_dma_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_dma_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (pixel_dma_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (pixel_dma_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (pixel_dma_avalon_pixel_source_data)                           //                        .data
	);

	gpu_qsys_pixel_fifo_mod pixel_fifo_mod (
		.clk_stream_in            (pll_outclk0_clk),                                      //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                       //         reset_stream_in.reset
		.clk_stream_out           (video_pll_vga_clk_clk),                                //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_001_reset_out_reset),                   //        reset_stream_out.reset
		.stream_in_ready          (pixel_dma_avalon_pixel_source_ready),                  //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (pixel_dma_avalon_pixel_source_startofpacket),          //                        .startofpacket
		.stream_in_endofpacket    (pixel_dma_avalon_pixel_source_endofpacket),            //                        .endofpacket
		.stream_in_valid          (pixel_dma_avalon_pixel_source_valid),                  //                        .valid
		.stream_in_data           (pixel_dma_avalon_pixel_source_data),                   //                        .data
		.stream_out_ready         (pixel_fifo_mod_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (pixel_fifo_mod_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (pixel_fifo_mod_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (pixel_fifo_mod_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (pixel_fifo_mod_avalon_dc_buffer_source_data)           //                        .data
	);

	gpu_qsys_pll pll (
		.refclk   (clk_clk),         //  refclk.clk
		.rst      (reset_reset),     //   reset.reset
		.outclk_0 (pll_outclk0_clk), // outclk0.clk
		.locked   ()                 // (terminated)
	);

	gpu_qsys_prim_assembly_fifo prim_assembly_fifo (
		.wrclock                       (pll_outclk0_clk),                                        //    clk_in.clk
		.wrreset_n                     (~rst_controller_reset_out_reset),                        //  reset_in.reset_n
		.rdclock                       (pll_outclk0_clk),                                        //   clk_out.clk
		.rdreset_n                     (~rst_controller_reset_out_reset),                        // reset_out.reset_n
		.avalonst_sink_valid           (prim_assembly_fifo_in_valid),                            //        in.valid
		.avalonst_sink_data            (prim_assembly_fifo_in_data),                             //          .data
		.avalonst_sink_ready           (prim_assembly_fifo_in_ready),                            //          .ready
		.avalonst_source_valid         (prim_assembly_fifo_out_valid),                           //       out.valid
		.avalonst_source_data          (prim_assembly_fifo_out_data),                            //          .data
		.avalonst_source_ready         (prim_assembly_fifo_out_ready),                           //          .ready
		.rdclk_control_slave_address   (mm_interconnect_2_prim_assembly_fifo_out_csr_address),   //   out_csr.address
		.rdclk_control_slave_read      (mm_interconnect_2_prim_assembly_fifo_out_csr_read),      //          .read
		.rdclk_control_slave_writedata (mm_interconnect_2_prim_assembly_fifo_out_csr_writedata), //          .writedata
		.rdclk_control_slave_write     (mm_interconnect_2_prim_assembly_fifo_out_csr_write),     //          .write
		.rdclk_control_slave_readdata  (mm_interconnect_2_prim_assembly_fifo_out_csr_readdata),  //          .readdata
		.wrclk_control_slave_address   (),                                                       //    in_csr.address
		.wrclk_control_slave_read      (),                                                       //          .read
		.wrclk_control_slave_writedata (),                                                       //          .writedata
		.wrclk_control_slave_write     (),                                                       //          .write
		.wrclk_control_slave_readdata  ()                                                        //          .readdata
	);

	gpu_qsys_prim_assembly_fifo raster_fifo (
		.wrclock                       (pll_outclk0_clk),                                 //    clk_in.clk
		.wrreset_n                     (~rst_controller_reset_out_reset),                 //  reset_in.reset_n
		.rdclock                       (pll_outclk0_clk),                                 //   clk_out.clk
		.rdreset_n                     (~rst_controller_reset_out_reset),                 // reset_out.reset_n
		.avalonst_sink_valid           (raster_fifo_in_valid),                            //        in.valid
		.avalonst_sink_data            (raster_fifo_in_data),                             //          .data
		.avalonst_sink_ready           (raster_fifo_in_ready),                            //          .ready
		.avalonst_source_valid         (raster_fifo_out_valid),                           //       out.valid
		.avalonst_source_data          (raster_fifo_out_data),                            //          .data
		.avalonst_source_ready         (raster_fifo_out_ready),                           //          .ready
		.rdclk_control_slave_address   (mm_interconnect_2_raster_fifo_out_csr_address),   //   out_csr.address
		.rdclk_control_slave_read      (mm_interconnect_2_raster_fifo_out_csr_read),      //          .read
		.rdclk_control_slave_writedata (mm_interconnect_2_raster_fifo_out_csr_writedata), //          .writedata
		.rdclk_control_slave_write     (mm_interconnect_2_raster_fifo_out_csr_write),     //          .write
		.rdclk_control_slave_readdata  (mm_interconnect_2_raster_fifo_out_csr_readdata),  //          .readdata
		.wrclk_control_slave_address   (),                                                //    in_csr.address
		.wrclk_control_slave_read      (),                                                //          .read
		.wrclk_control_slave_writedata (),                                                //          .writedata
		.wrclk_control_slave_write     (),                                                //          .write
		.wrclk_control_slave_readdata  ()                                                 //          .readdata
	);

	gpu_qsys_prim_assembly_fifo vert_processing_fifo (
		.wrclock                       (pll_outclk0_clk),                                          //    clk_in.clk
		.wrreset_n                     (~rst_controller_reset_out_reset),                          //  reset_in.reset_n
		.rdclock                       (pll_outclk0_clk),                                          //   clk_out.clk
		.rdreset_n                     (~rst_controller_reset_out_reset),                          // reset_out.reset_n
		.avalonst_sink_valid           (vert_processing_fifo_in_valid),                            //        in.valid
		.avalonst_sink_data            (vert_processing_fifo_in_data),                             //          .data
		.avalonst_sink_ready           (vert_processing_fifo_in_ready),                            //          .ready
		.avalonst_source_valid         (vert_processing_fifo_out_valid),                           //       out.valid
		.avalonst_source_data          (vert_processing_fifo_out_data),                            //          .data
		.avalonst_source_ready         (vert_processing_fifo_out_ready),                           //          .ready
		.rdclk_control_slave_address   (mm_interconnect_2_vert_processing_fifo_out_csr_address),   //   out_csr.address
		.rdclk_control_slave_read      (mm_interconnect_2_vert_processing_fifo_out_csr_read),      //          .read
		.rdclk_control_slave_writedata (mm_interconnect_2_vert_processing_fifo_out_csr_writedata), //          .writedata
		.rdclk_control_slave_write     (mm_interconnect_2_vert_processing_fifo_out_csr_write),     //          .write
		.rdclk_control_slave_readdata  (mm_interconnect_2_vert_processing_fifo_out_csr_readdata),  //          .readdata
		.wrclk_control_slave_address   (),                                                         //    in_csr.address
		.wrclk_control_slave_read      (),                                                         //          .read
		.wrclk_control_slave_writedata (),                                                         //          .writedata
		.wrclk_control_slave_write     (),                                                         //          .write
		.wrclk_control_slave_readdata  ()                                                          //          .readdata
	);

	gpu_qsys_vga_controller vga_controller (
		.clk           (video_pll_vga_clk_clk),                                //                clk.clk
		.reset         (rst_controller_001_reset_out_reset),                   //              reset.reset
		.data          (pixel_fifo_mod_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (pixel_fifo_mod_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (pixel_fifo_mod_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (pixel_fifo_mod_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (pixel_fifo_mod_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_controller_external_interface_CLK),                // external_interface.export
		.VGA_HS        (vga_controller_external_interface_HS),                 //                   .export
		.VGA_VS        (vga_controller_external_interface_VS),                 //                   .export
		.VGA_BLANK     (vga_controller_external_interface_BLANK),              //                   .export
		.VGA_SYNC      (vga_controller_external_interface_SYNC),               //                   .export
		.VGA_R         (vga_controller_external_interface_R),                  //                   .export
		.VGA_G         (vga_controller_external_interface_G),                  //                   .export
		.VGA_B         (vga_controller_external_interface_B)                   //                   .export
	);

	gpu_qsys_video_pll video_pll (
		.ref_clk_clk        (video_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (~hps_h2f_reset_reset),         //    ref_reset.reset
		.vga_clk_clk        (video_pll_vga_clk_clk),        //      vga_clk.clk
		.reset_source_reset (video_pll_reset_source_reset)  // reset_source.reset
	);

	gpu_qsys_mm_interconnect_0 mm_interconnect_0 (
		.pll_outclk0_clk                                    (pll_outclk0_clk),                                                      //                          pll_outclk0.clk
		.gpu_main_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                                       // gpu_main_reset_reset_bridge_in_reset.reset
		.gpu_main_avalon_master_address                     (gpu_main_avalon_master_address),                                       //               gpu_main_avalon_master.address
		.gpu_main_avalon_master_waitrequest                 (gpu_main_avalon_master_waitrequest),                                   //                                     .waitrequest
		.gpu_main_avalon_master_byteenable                  (gpu_main_avalon_master_byteenable),                                    //                                     .byteenable
		.gpu_main_avalon_master_read                        (gpu_main_avalon_master_read),                                          //                                     .read
		.gpu_main_avalon_master_readdata                    (gpu_main_avalon_master_readdata),                                      //                                     .readdata
		.gpu_main_avalon_master_write                       (gpu_main_avalon_master_write),                                         //                                     .write
		.gpu_main_avalon_master_writedata                   (gpu_main_avalon_master_writedata),                                     //                                     .writedata
		.address_span_extender_windowed_slave_address       (mm_interconnect_0_address_span_extender_windowed_slave_address),       // address_span_extender_windowed_slave.address
		.address_span_extender_windowed_slave_write         (mm_interconnect_0_address_span_extender_windowed_slave_write),         //                                     .write
		.address_span_extender_windowed_slave_read          (mm_interconnect_0_address_span_extender_windowed_slave_read),          //                                     .read
		.address_span_extender_windowed_slave_readdata      (mm_interconnect_0_address_span_extender_windowed_slave_readdata),      //                                     .readdata
		.address_span_extender_windowed_slave_writedata     (mm_interconnect_0_address_span_extender_windowed_slave_writedata),     //                                     .writedata
		.address_span_extender_windowed_slave_burstcount    (mm_interconnect_0_address_span_extender_windowed_slave_burstcount),    //                                     .burstcount
		.address_span_extender_windowed_slave_byteenable    (mm_interconnect_0_address_span_extender_windowed_slave_byteenable),    //                                     .byteenable
		.address_span_extender_windowed_slave_readdatavalid (mm_interconnect_0_address_span_extender_windowed_slave_readdatavalid), //                                     .readdatavalid
		.address_span_extender_windowed_slave_waitrequest   (mm_interconnect_0_address_span_extender_windowed_slave_waitrequest)    //                                     .waitrequest
	);

	gpu_qsys_mm_interconnect_1 mm_interconnect_1 (
		.hps_f2h_axi_slave_awid                              (mm_interconnect_1_hps_f2h_axi_slave_awid),            //                     hps_f2h_axi_slave.awid
		.hps_f2h_axi_slave_awaddr                            (mm_interconnect_1_hps_f2h_axi_slave_awaddr),          //                                      .awaddr
		.hps_f2h_axi_slave_awlen                             (mm_interconnect_1_hps_f2h_axi_slave_awlen),           //                                      .awlen
		.hps_f2h_axi_slave_awsize                            (mm_interconnect_1_hps_f2h_axi_slave_awsize),          //                                      .awsize
		.hps_f2h_axi_slave_awburst                           (mm_interconnect_1_hps_f2h_axi_slave_awburst),         //                                      .awburst
		.hps_f2h_axi_slave_awlock                            (mm_interconnect_1_hps_f2h_axi_slave_awlock),          //                                      .awlock
		.hps_f2h_axi_slave_awcache                           (mm_interconnect_1_hps_f2h_axi_slave_awcache),         //                                      .awcache
		.hps_f2h_axi_slave_awprot                            (mm_interconnect_1_hps_f2h_axi_slave_awprot),          //                                      .awprot
		.hps_f2h_axi_slave_awuser                            (mm_interconnect_1_hps_f2h_axi_slave_awuser),          //                                      .awuser
		.hps_f2h_axi_slave_awvalid                           (mm_interconnect_1_hps_f2h_axi_slave_awvalid),         //                                      .awvalid
		.hps_f2h_axi_slave_awready                           (mm_interconnect_1_hps_f2h_axi_slave_awready),         //                                      .awready
		.hps_f2h_axi_slave_wid                               (mm_interconnect_1_hps_f2h_axi_slave_wid),             //                                      .wid
		.hps_f2h_axi_slave_wdata                             (mm_interconnect_1_hps_f2h_axi_slave_wdata),           //                                      .wdata
		.hps_f2h_axi_slave_wstrb                             (mm_interconnect_1_hps_f2h_axi_slave_wstrb),           //                                      .wstrb
		.hps_f2h_axi_slave_wlast                             (mm_interconnect_1_hps_f2h_axi_slave_wlast),           //                                      .wlast
		.hps_f2h_axi_slave_wvalid                            (mm_interconnect_1_hps_f2h_axi_slave_wvalid),          //                                      .wvalid
		.hps_f2h_axi_slave_wready                            (mm_interconnect_1_hps_f2h_axi_slave_wready),          //                                      .wready
		.hps_f2h_axi_slave_bid                               (mm_interconnect_1_hps_f2h_axi_slave_bid),             //                                      .bid
		.hps_f2h_axi_slave_bresp                             (mm_interconnect_1_hps_f2h_axi_slave_bresp),           //                                      .bresp
		.hps_f2h_axi_slave_bvalid                            (mm_interconnect_1_hps_f2h_axi_slave_bvalid),          //                                      .bvalid
		.hps_f2h_axi_slave_bready                            (mm_interconnect_1_hps_f2h_axi_slave_bready),          //                                      .bready
		.hps_f2h_axi_slave_arid                              (mm_interconnect_1_hps_f2h_axi_slave_arid),            //                                      .arid
		.hps_f2h_axi_slave_araddr                            (mm_interconnect_1_hps_f2h_axi_slave_araddr),          //                                      .araddr
		.hps_f2h_axi_slave_arlen                             (mm_interconnect_1_hps_f2h_axi_slave_arlen),           //                                      .arlen
		.hps_f2h_axi_slave_arsize                            (mm_interconnect_1_hps_f2h_axi_slave_arsize),          //                                      .arsize
		.hps_f2h_axi_slave_arburst                           (mm_interconnect_1_hps_f2h_axi_slave_arburst),         //                                      .arburst
		.hps_f2h_axi_slave_arlock                            (mm_interconnect_1_hps_f2h_axi_slave_arlock),          //                                      .arlock
		.hps_f2h_axi_slave_arcache                           (mm_interconnect_1_hps_f2h_axi_slave_arcache),         //                                      .arcache
		.hps_f2h_axi_slave_arprot                            (mm_interconnect_1_hps_f2h_axi_slave_arprot),          //                                      .arprot
		.hps_f2h_axi_slave_aruser                            (mm_interconnect_1_hps_f2h_axi_slave_aruser),          //                                      .aruser
		.hps_f2h_axi_slave_arvalid                           (mm_interconnect_1_hps_f2h_axi_slave_arvalid),         //                                      .arvalid
		.hps_f2h_axi_slave_arready                           (mm_interconnect_1_hps_f2h_axi_slave_arready),         //                                      .arready
		.hps_f2h_axi_slave_rid                               (mm_interconnect_1_hps_f2h_axi_slave_rid),             //                                      .rid
		.hps_f2h_axi_slave_rdata                             (mm_interconnect_1_hps_f2h_axi_slave_rdata),           //                                      .rdata
		.hps_f2h_axi_slave_rresp                             (mm_interconnect_1_hps_f2h_axi_slave_rresp),           //                                      .rresp
		.hps_f2h_axi_slave_rlast                             (mm_interconnect_1_hps_f2h_axi_slave_rlast),           //                                      .rlast
		.hps_f2h_axi_slave_rvalid                            (mm_interconnect_1_hps_f2h_axi_slave_rvalid),          //                                      .rvalid
		.hps_f2h_axi_slave_rready                            (mm_interconnect_1_hps_f2h_axi_slave_rready),          //                                      .rready
		.pll_outclk0_clk                                     (pll_outclk0_clk),                                     //                           pll_outclk0.clk
		.pixel_dma_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                      // pixel_dma_reset_reset_bridge_in_reset.reset
		.address_span_extender_expanded_master_address       (address_span_extender_expanded_master_address),       // address_span_extender_expanded_master.address
		.address_span_extender_expanded_master_waitrequest   (address_span_extender_expanded_master_waitrequest),   //                                      .waitrequest
		.address_span_extender_expanded_master_burstcount    (address_span_extender_expanded_master_burstcount),    //                                      .burstcount
		.address_span_extender_expanded_master_byteenable    (address_span_extender_expanded_master_byteenable),    //                                      .byteenable
		.address_span_extender_expanded_master_read          (address_span_extender_expanded_master_read),          //                                      .read
		.address_span_extender_expanded_master_readdata      (address_span_extender_expanded_master_readdata),      //                                      .readdata
		.address_span_extender_expanded_master_readdatavalid (address_span_extender_expanded_master_readdatavalid), //                                      .readdatavalid
		.address_span_extender_expanded_master_write         (address_span_extender_expanded_master_write),         //                                      .write
		.address_span_extender_expanded_master_writedata     (address_span_extender_expanded_master_writedata),     //                                      .writedata
		.pixel_dma_avalon_pixel_dma_master_address           (pixel_dma_avalon_pixel_dma_master_address),           //     pixel_dma_avalon_pixel_dma_master.address
		.pixel_dma_avalon_pixel_dma_master_waitrequest       (pixel_dma_avalon_pixel_dma_master_waitrequest),       //                                      .waitrequest
		.pixel_dma_avalon_pixel_dma_master_read              (pixel_dma_avalon_pixel_dma_master_read),              //                                      .read
		.pixel_dma_avalon_pixel_dma_master_readdata          (pixel_dma_avalon_pixel_dma_master_readdata),          //                                      .readdata
		.pixel_dma_avalon_pixel_dma_master_readdatavalid     (pixel_dma_avalon_pixel_dma_master_readdatavalid),     //                                      .readdatavalid
		.pixel_dma_avalon_pixel_dma_master_lock              (pixel_dma_avalon_pixel_dma_master_lock)               //                                      .lock
	);

	gpu_qsys_mm_interconnect_2 mm_interconnect_2 (
		.hps_h2f_axi_master_awid                     (hps_h2f_axi_master_awid),                                     //                    hps_h2f_axi_master.awid
		.hps_h2f_axi_master_awaddr                   (hps_h2f_axi_master_awaddr),                                   //                                      .awaddr
		.hps_h2f_axi_master_awlen                    (hps_h2f_axi_master_awlen),                                    //                                      .awlen
		.hps_h2f_axi_master_awsize                   (hps_h2f_axi_master_awsize),                                   //                                      .awsize
		.hps_h2f_axi_master_awburst                  (hps_h2f_axi_master_awburst),                                  //                                      .awburst
		.hps_h2f_axi_master_awlock                   (hps_h2f_axi_master_awlock),                                   //                                      .awlock
		.hps_h2f_axi_master_awcache                  (hps_h2f_axi_master_awcache),                                  //                                      .awcache
		.hps_h2f_axi_master_awprot                   (hps_h2f_axi_master_awprot),                                   //                                      .awprot
		.hps_h2f_axi_master_awvalid                  (hps_h2f_axi_master_awvalid),                                  //                                      .awvalid
		.hps_h2f_axi_master_awready                  (hps_h2f_axi_master_awready),                                  //                                      .awready
		.hps_h2f_axi_master_wid                      (hps_h2f_axi_master_wid),                                      //                                      .wid
		.hps_h2f_axi_master_wdata                    (hps_h2f_axi_master_wdata),                                    //                                      .wdata
		.hps_h2f_axi_master_wstrb                    (hps_h2f_axi_master_wstrb),                                    //                                      .wstrb
		.hps_h2f_axi_master_wlast                    (hps_h2f_axi_master_wlast),                                    //                                      .wlast
		.hps_h2f_axi_master_wvalid                   (hps_h2f_axi_master_wvalid),                                   //                                      .wvalid
		.hps_h2f_axi_master_wready                   (hps_h2f_axi_master_wready),                                   //                                      .wready
		.hps_h2f_axi_master_bid                      (hps_h2f_axi_master_bid),                                      //                                      .bid
		.hps_h2f_axi_master_bresp                    (hps_h2f_axi_master_bresp),                                    //                                      .bresp
		.hps_h2f_axi_master_bvalid                   (hps_h2f_axi_master_bvalid),                                   //                                      .bvalid
		.hps_h2f_axi_master_bready                   (hps_h2f_axi_master_bready),                                   //                                      .bready
		.hps_h2f_axi_master_arid                     (hps_h2f_axi_master_arid),                                     //                                      .arid
		.hps_h2f_axi_master_araddr                   (hps_h2f_axi_master_araddr),                                   //                                      .araddr
		.hps_h2f_axi_master_arlen                    (hps_h2f_axi_master_arlen),                                    //                                      .arlen
		.hps_h2f_axi_master_arsize                   (hps_h2f_axi_master_arsize),                                   //                                      .arsize
		.hps_h2f_axi_master_arburst                  (hps_h2f_axi_master_arburst),                                  //                                      .arburst
		.hps_h2f_axi_master_arlock                   (hps_h2f_axi_master_arlock),                                   //                                      .arlock
		.hps_h2f_axi_master_arcache                  (hps_h2f_axi_master_arcache),                                  //                                      .arcache
		.hps_h2f_axi_master_arprot                   (hps_h2f_axi_master_arprot),                                   //                                      .arprot
		.hps_h2f_axi_master_arvalid                  (hps_h2f_axi_master_arvalid),                                  //                                      .arvalid
		.hps_h2f_axi_master_arready                  (hps_h2f_axi_master_arready),                                  //                                      .arready
		.hps_h2f_axi_master_rid                      (hps_h2f_axi_master_rid),                                      //                                      .rid
		.hps_h2f_axi_master_rdata                    (hps_h2f_axi_master_rdata),                                    //                                      .rdata
		.hps_h2f_axi_master_rresp                    (hps_h2f_axi_master_rresp),                                    //                                      .rresp
		.hps_h2f_axi_master_rlast                    (hps_h2f_axi_master_rlast),                                    //                                      .rlast
		.hps_h2f_axi_master_rvalid                   (hps_h2f_axi_master_rvalid),                                   //                                      .rvalid
		.hps_h2f_axi_master_rready                   (hps_h2f_axi_master_rready),                                   //                                      .rready
		.pll_outclk0_clk                             (pll_outclk0_clk),                                             //                           pll_outclk0.clk
		.pixel_dma_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // pixel_dma_reset_reset_bridge_in_reset.reset
		.instr_fifo_in_address                       (mm_interconnect_2_instr_fifo_in_address),                     //                         instr_fifo_in.address
		.instr_fifo_in_write                         (mm_interconnect_2_instr_fifo_in_write),                       //                                      .write
		.instr_fifo_in_writedata                     (mm_interconnect_2_instr_fifo_in_writedata),                   //                                      .writedata
		.instr_fifo_in_waitrequest                   (mm_interconnect_2_instr_fifo_in_waitrequest),                 //                                      .waitrequest
		.instr_fifo_in_csr_address                   (mm_interconnect_2_instr_fifo_in_csr_address),                 //                     instr_fifo_in_csr.address
		.instr_fifo_in_csr_write                     (mm_interconnect_2_instr_fifo_in_csr_write),                   //                                      .write
		.instr_fifo_in_csr_read                      (mm_interconnect_2_instr_fifo_in_csr_read),                    //                                      .read
		.instr_fifo_in_csr_readdata                  (mm_interconnect_2_instr_fifo_in_csr_readdata),                //                                      .readdata
		.instr_fifo_in_csr_writedata                 (mm_interconnect_2_instr_fifo_in_csr_writedata),               //                                      .writedata
		.pixel_dma_avalon_control_slave_address      (mm_interconnect_2_pixel_dma_avalon_control_slave_address),    //        pixel_dma_avalon_control_slave.address
		.pixel_dma_avalon_control_slave_write        (mm_interconnect_2_pixel_dma_avalon_control_slave_write),      //                                      .write
		.pixel_dma_avalon_control_slave_read         (mm_interconnect_2_pixel_dma_avalon_control_slave_read),       //                                      .read
		.pixel_dma_avalon_control_slave_readdata     (mm_interconnect_2_pixel_dma_avalon_control_slave_readdata),   //                                      .readdata
		.pixel_dma_avalon_control_slave_writedata    (mm_interconnect_2_pixel_dma_avalon_control_slave_writedata),  //                                      .writedata
		.pixel_dma_avalon_control_slave_byteenable   (mm_interconnect_2_pixel_dma_avalon_control_slave_byteenable), //                                      .byteenable
		.prim_assembly_fifo_out_csr_address          (mm_interconnect_2_prim_assembly_fifo_out_csr_address),        //            prim_assembly_fifo_out_csr.address
		.prim_assembly_fifo_out_csr_write            (mm_interconnect_2_prim_assembly_fifo_out_csr_write),          //                                      .write
		.prim_assembly_fifo_out_csr_read             (mm_interconnect_2_prim_assembly_fifo_out_csr_read),           //                                      .read
		.prim_assembly_fifo_out_csr_readdata         (mm_interconnect_2_prim_assembly_fifo_out_csr_readdata),       //                                      .readdata
		.prim_assembly_fifo_out_csr_writedata        (mm_interconnect_2_prim_assembly_fifo_out_csr_writedata),      //                                      .writedata
		.raster_fifo_out_csr_address                 (mm_interconnect_2_raster_fifo_out_csr_address),               //                   raster_fifo_out_csr.address
		.raster_fifo_out_csr_write                   (mm_interconnect_2_raster_fifo_out_csr_write),                 //                                      .write
		.raster_fifo_out_csr_read                    (mm_interconnect_2_raster_fifo_out_csr_read),                  //                                      .read
		.raster_fifo_out_csr_readdata                (mm_interconnect_2_raster_fifo_out_csr_readdata),              //                                      .readdata
		.raster_fifo_out_csr_writedata               (mm_interconnect_2_raster_fifo_out_csr_writedata),             //                                      .writedata
		.vert_processing_fifo_out_csr_address        (mm_interconnect_2_vert_processing_fifo_out_csr_address),      //          vert_processing_fifo_out_csr.address
		.vert_processing_fifo_out_csr_write          (mm_interconnect_2_vert_processing_fifo_out_csr_write),        //                                      .write
		.vert_processing_fifo_out_csr_read           (mm_interconnect_2_vert_processing_fifo_out_csr_read),         //                                      .read
		.vert_processing_fifo_out_csr_readdata       (mm_interconnect_2_vert_processing_fifo_out_csr_readdata),     //                                      .readdata
		.vert_processing_fifo_out_csr_writedata      (mm_interconnect_2_vert_processing_fifo_out_csr_writedata)     //                                      .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_h2f_reset_reset),           // reset_in0.reset
		.clk            (pll_outclk0_clk),                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_h2f_reset_reset),               // reset_in0.reset
		.reset_in1      (video_pll_reset_source_reset),       // reset_in1.reset
		.clk            (video_pll_vga_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
